module pipeline();

endmodule;